module decoder
(
    input clk,
    input wire [7:0] instr,
    output reg [1:0] alu_op1_sel,
    output reg [1:0] alu_op2_sel,
);

    always @(posedge clk) begin

    end

endmodule

module regfile
(
    input wire clk,
    output reg [7:0] acc_reg,
    output reg [7:0] x_reg,
    output reg [7:0] y_reg,
    output reg [15:0] pc,
    output reg [7:0] status_reg
);

    always @(posedge clk) begin
        pc <= pc + 1;
    end

endmodule

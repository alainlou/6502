module regfile
(

)

endmodule regfile

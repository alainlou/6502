`ifndef TYPES_GUARD_DEF
`define TYPES_GUARD_DEF

package types;
    typedef enum bit [1:0] { X_REG, Y_REG, ACC_REG } reg_t;
endpackage

`endif

module code_mem #
(
    param NUM_BYTES=1024
)
(
    input wire [15:0] rdaddr,
    output wire []
)

module top
(
    input FPGA_CLK,
    input UART_RXD,
    output UART_TXD
);



endmodule
